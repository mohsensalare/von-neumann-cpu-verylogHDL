`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:25:52 11/02/2020 
// Design Name: 
// Module Name:    SC_M 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module SC_M(
    input clk,
    input rst,
    input rstsc,
    output [2:0] DATA_out
    );
	reg counter[2:0];

endmodule
